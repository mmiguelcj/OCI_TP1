library verilog;
use verilog.vl_types.all;
entity KronosX is
    port(
        pin_name5       : out    vl_logic;
        pin_name1       : in     vl_logic;
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic
    );
end KronosX;
