library verilog;
use verilog.vl_types.all;
entity KronosX_vlg_check_tst is
    port(
        pin_name5       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end KronosX_vlg_check_tst;
