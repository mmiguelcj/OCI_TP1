library verilog;
use verilog.vl_types.all;
entity Shift_vlg_vec_tst is
end Shift_vlg_vec_tst;
