library verilog;
use verilog.vl_types.all;
entity KronosX_vlg_vec_tst is
end KronosX_vlg_vec_tst;
